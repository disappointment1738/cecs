
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: CSULB
// Engineer: Amin Rezaei
// Create Date: 08/22/2020 06:59:39 PM
// Design Name: 361_Lab1
// Module Name: ArrMult_4bit
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module ArrMult_4bit(
  input [3:0] a, b,
  output [7:0] prod
  );
    wire [10:0] carry;
    wire [5:0] partialSum;

    //Partial Products
    wire [3:0] pp [0:3];

    //Asign Patrial Products
    //row 0
    mux2to1 m00(.a(a[0]), .b(1'b0), .sel(b[0]), .out(pp[0][0]));
    mux2to1 m01(.a(a[1]), .b(1'b0), .sel(b[0]), .out(pp[0][1]));
    mux2to1 m02(.a(a[2]), .b(1'b0), .sel(b[0]), .out(pp[0][2]));
    mux2to1 m03(.a(a[3]), .b(1'b0), .sel(b[0]), .out(pp[0][3]));
    //row 1
    //row 2
    //row 3

    //Assign Adding Circuit
    //sum 0
    assign prod[0] = pp[0][0];
    //sum 1
    HA h0(.a(pp[1][0]), .b(pp[0][1]), .c_out(carry[0]), .sum(prod[1]));
    //sum 2
    FA f0(.a(pp[1][1]), .b(pp[0][2]), .c_in(carry[0]), .c_out(carry[1]), .sum(partialSum[0]));
    HA h1(.a(pp[2][0]), .b(partialSum[0]), .c_out(carry[2]), .sum(prod[2]));
    //sum 3
    //sum 4
    //sum 5
    //sum 6 & sum 7
    
endmodule
